`timescale 1ns / 1ps

// this adapts the clock module to the main state machine

module clock_main_adp(clk,rst,en,toggle_btn);
endmodule
